library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity instruction_memory is
  port (
    address     : in    std_logic_vector(31 downto 0);
    instruction : out   std_logic_vector(31 downto 0)
  );
end entity instruction_memory;

architecture behavioral of instruction_memory is

  type instruction_array is array (0 to 127) of std_logic_vector(31 downto 0);

  signal instructions : instruction_array := (
0 => "00000000000000000000000000000000",
 1 => "00000000000000000000000000000000",
 2 => "00100000000010000000000000000000",
 3 => "10101111101010000000000000000000",
 4 => "00100000000010000000000000000001",
 5 => "10101111101010000000000000000100",
 6 => "00100000000010000000000000000001",
 7 => "10101111101010000000000000001000",
 8 => "00100000000010000000000000000010",
 9 => "10101111101010000000000000001100",
10 => "00100000000010000000000000000011",
11 => "10101111101010000000000000010000",
12 => "00100000000010000000000000000101",
13 => "10101111101010000000000000010100",
14 => "00100000000010000000000000001000",
15 => "10101111101010000000000000011000",
16 => "00100000000010000000000000001101",
17 => "10101111101010000000000000011100",
18 => "00100000000010000000000000010101",
19 => "10101111101010000000000000100000",
20 => "00100000000010000000000000100010",
21 => "10101111101010000000000000100100",
22 => "00100000000010000000000000110111",
23 => "10101111101010000000000000101000",
24 => "00100000000010000000000001011001",
25 => "10101111101010000000000000101100",
26 => "00100000000010000000000010010000",
27 => "10101111101010000000000000110000",
28 => "00100000000010000000000011101001",
29 => "10101111101010000000000000110100",
30 => "00100000000010000000000101111001",
31 => "10101111101010000000000000111000",
32 => "00100000000010000000001001100010",
33 => "10101111101010000000000000111100",
34=>  "00001000000000000000000000100010",
35 to 127=> (others => '0'));

begin

  instruction <= instructions(to_integer(unsigned(address(31 downto 2))));

end architecture behavioral;
